-- Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, the Altera Quartus Prime License Agreement,
-- the Altera MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Altera and sold by Altera or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- Generated by Quartus Prime Version 16.0.0 Build 211 04/27/2016 SJ Lite Edition
-- Created on Tue Sep 25 08:46:49 2018

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY fsm_relogio IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        US_MAX : IN STD_LOGIC := '0';
        DS_GO : IN STD_LOGIC := '0';
        DS_MAX : IN STD_LOGIC := '0';
        UM_GO : IN STD_LOGIC := '0';
        UM_MAX : IN STD_LOGIC := '0';
        DM_GO : IN STD_LOGIC := '0';
        DM_MAX : IN STD_LOGIC := '0';
        UH_GO : IN STD_LOGIC := '0';
        UH_MAX : IN STD_LOGIC := '0';
        DH_GO : IN STD_LOGIC := '0';
        DH_MAX : IN STD_LOGIC := '0';
        Clock_Restart : IN STD_LOGIC := '0';
        palavra : OUT STD_LOGIC_VECTOR(12 DOWNTO 0)
    );
END fsm_relogio;

ARCHITECTURE BEHAVIOR OF fsm_relogio IS
    TYPE type_fstate IS (conta_segundo,Incrementa_DS_parte_I,incrementa_DS_parteII,zera_DS,conta_minuto,incrementa_DM_parte_I,incrementa_DM_parte_II,zera_DM,conta_hora,incrementa_DH_parte_I,incrementa_DH_parte_II,zera_DH);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,US_MAX,DS_GO,DS_MAX,UM_GO,UM_MAX,DM_GO,DM_MAX,UH_GO,UH_MAX,DH_GO,DH_MAX,Clock_Restart)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= conta_segundo;
            palavra <= "0000000000000";
        ELSE
            palavra <= "0000000000000";
            CASE fstate IS
                WHEN conta_segundo =>
                    IF ((US_MAX = '1')) THEN
                        reg_fstate <= Incrementa_DS_parte_I;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= conta_segundo;
                    END IF;

                    palavra <= "0000000110000";
                WHEN Incrementa_DS_parte_I =>
                    reg_fstate <= incrementa_DS_parteII;

                    palavra <= "0010000101000";
                WHEN incrementa_DS_parteII =>
                    IF ((DS_MAX = '1')) THEN
                        reg_fstate <= zera_DS;
                    ELSIF (NOT((DS_MAX = '1'))) THEN
                        reg_fstate <= conta_segundo;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= incrementa_DS_parteII;
                    END IF;

                    palavra <= "0000001000001";
                WHEN zera_DS =>
                    reg_fstate <= conta_minuto;

                    palavra <= "0010001011001";
                WHEN conta_minuto =>
                    IF ((UM_MAX = '1')) THEN
                        reg_fstate <= incrementa_DM_parte_I;
                    ELSIF (NOT((UM_MAX = '1'))) THEN
                        reg_fstate <= conta_segundo;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= conta_minuto;
                    END IF;

                    palavra <= "0000010000010";
                WHEN incrementa_DM_parte_I =>
                    reg_fstate <= incrementa_DM_parte_II;

                    palavra <= "0010010101010";
                WHEN incrementa_DM_parte_II =>
                    IF ((DM_MAX = '1')) THEN
                        reg_fstate <= zera_DM;
                    ELSIF (NOT((DM_MAX = '1'))) THEN
                        reg_fstate <= conta_minuto;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= incrementa_DM_parte_II;
                    END IF;

                    palavra <= "0000011000011";
                WHEN zera_DM =>
                    reg_fstate <= conta_hora;

                    palavra <= "0010011011011";
                WHEN conta_hora =>
                    IF ((UH_MAX = '1')) THEN
                        reg_fstate <= incrementa_DH_parte_I;
                    ELSIF (NOT((UH_MAX = '1'))) THEN
                        reg_fstate <= conta_segundo;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= conta_hora;
                    END IF;

                    palavra <= "0000100000100";
                WHEN incrementa_DH_parte_I =>
                    reg_fstate <= incrementa_DH_parte_II;

                    palavra <= "0010100001100";
                WHEN incrementa_DH_parte_II =>
                    IF ((DH_MAX = '1')) THEN
                        reg_fstate <= zera_DH;
                    ELSIF (NOT((DH_MAX = '1'))) THEN
                        reg_fstate <= conta_hora;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= incrementa_DH_parte_II;
                    END IF;
						  
						  palavra <= "0000101000101";
                WHEN zera_DH =>
                    IF ((Clock_Restart = '1')) THEN
                        reg_fstate <= conta_segundo;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= zera_DH;
                    END IF;

                    palavra <= "0010101010101";
                WHEN OTHERS => 
                    palavra <= "XXXXXXXXXXXXX";
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
